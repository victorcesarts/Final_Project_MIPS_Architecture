library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all; 

entity InstrMemory is 
    port(
        address : in std_logic_vector(31 downto 0);
        instr : out std_logic_vector(31 downto 0)
    );
end InstrMemory;
--addi $16,$16,0x0000000       	
--add $4,$16,$0            	
--jal 0x0040001c           	
--add $17,$2,$0            	
--addiu $2,$0,0x0000000a   
--syscall                  
--addi $29,$29,0xfffffff   
--sw $8,0x0000000c($29)    
--sw $9,0x00000008($29)    
--sw $10,0x00000004($29)   
--sw $11,0x00000000($29)   
--addi $8,$0,0x00000001    
--slt $9,$8,$4             
--beq $9,$0,0x00000008     	
--add $10,$4,$0            		
--add $11,$8,$0            	
--slt $9,$8,$10            	
--beq $9,$0,0x00000007     	
--mult $11,$8              	
--mflo $11                 	
--addi $8,$8,0x00000001    	
--j 0x00400044             	
--addi $11,$0,0x00000001   	
--addu $2,$0,$11           	
--j 0x00400078             	
--mult $11,$4              	
--mflo $11                 	
--addu $2,$0,$11           	
--j 0x00400078             	
--lw $8,0x0000000c($29)    	
--lw $9,0x00000008($29)    	
--lw $10,0x00000004($29)   	
--lw $11,0x00000000($29)   	
--addi $29,$29,0x0000001   	
--jr $31 

architecture InstrARCH of InstrMemory is 
signal rom_addr : std_logic_vector(7 downto 0);
type rom is array (0 to 34) of std_logic_vector(31 downto 0);

constant Instr_data : 
rom :=rom'(
"00100010000100000000000000001100",
"00000010000000000010000000100000",
"00001100000100000000000000000111",
"00000000010000001000100000100000",
"00100100000000100000000000001010",
"00000000000000000000000000001100",
"00100011101111011111111111110000",
"10101111101010000000000000001100",
"10101111101010010000000000001000",
"10101111101010100000000000000100",
"10101111101010110000000000000000",
"00100000000010000000000000000001",
"00000001000001000100100000101010",
"00010001001000000000000000001000",
"00000000100000000101000000100000",
"00000001000000000101100000100000",
"00000001000010100100100000101010",
"00010001001000000000000000000111",
"00000001011010000000000000011000",
"00000000000000000101100000010010",
"00100001000010000000000000000001",
"00001000000100000000000000010001",
"00100000000010110000000000000001",
"00000000000010110001000000100001",
"00001000000100000000000000011110",
"00000001011001000000000000011000",
"00000000000000000101100000010010",
"00000000000010110001000000100001",
"00001000000100000000000000011110",
"10001111101010000000000000001100",
"10001111101010010000000000001000",
"10001111101010100000000000000100",
"10001111101010110000000000000000",
"00100011101111010000000000010000",
"00000011111000000000000000001000");
begin
    rom_addr <= address(9 downto 2);
    instr <= Instr_data(to_integer(unsigned(rom_addr))) when ((address >= x"00400000") and (address <= x"0FFFFFFD")) else x"00000000";      
end InstrARCH; 